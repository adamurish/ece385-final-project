module AppleIIe ;