module AppleIIe ();